package decode_test_pkg;
 
	import uvm_pkg::*;
        import uvmf_base_pkg::*;
	`include "uvm_macros.svh"
	import decode_env_pkg::*;
	import decode_in_pkg::*;
	import decode_out_pkg::*;
		
	`include "decode_test_pkg/print_component.sv"
	 `include "decode_test_pkg/test_top.svh"
	
	
endpackage
